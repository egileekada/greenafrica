<svg 
xmlns="http://www.w3.org/2000/svg" 
width="10.828" height="6.414" 
viewBox="0 0 10.828 6.414">
<defs>
</defs>
<path 
 fill="none"
 stroke-linecap="round"
 stroke-linejoin="round"
 stroke-width="2px"
 d="M864.559,93l4,4,4-4" 
 transform="translate(-863.145 -91.586)"/>
</svg>